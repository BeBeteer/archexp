`timescale 1ns / 1ps

module Alu (
		input [31:0] inputA,
		input [31:0] inputB,
		input [3:0] operation,
		output [31:0] output_
	);

	assign output_ =
			operation == ALU_ADD ? $signed(inputA) + $signed(inputB)
			: operation == ALU_ADDU ? inputA + inputB
			: operation == ALU_SUB ? $signed(inputA) - $signed(inputB)
			: operation == ALU_SUBU ? inputA - inputB
			: operation == ALU_AND ? inputA & inputB
			: operation == ALU_OR ? inputA | inputB
			: operation == ALU_XOR ? inputA ^ inputB
			: operation == ALU_NOR ? ~(inputA | inputB)
			: operation == ALU_SLL ? inputB << inputA
			: operation == ALU_SRL ? inputB >> inputA
			: operation == ALU_SRA ? inputB >>> inputA
			: 32'b0;
endmodule
